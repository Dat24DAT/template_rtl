module #{DESIGN_NAME} (
   
);
  
endmodule
