
module #{DESIGN_NAME}_tb;

// Parameters
localparam integer CLK_PERIOD = 10000;
//Declare Ports

//instantiate DUT here

////

always #(CLK_PERIOD / 2) clk = !clk;
initial begin
  intialize_input_values();
  reset();
  //give inputs at the negedge of the clock here
  @(negedge clk);
 
  $finish();
end
////utility tasks
task reset();
  rst_n = 0;
  #(3 * CLK_PERIOD);
  rst_n = 1;
  @(negedge clk);
endtask

task intialize_input_values();
  clk = 0;
  // all inputs to zero here
  en  = 1'b0;
endtask

task check_outputs(input logic [0:2] outputs, input logic [0:2] expected_outputs);
  @(negedge clk);
  assert (outputs === expected_outputs) begin
    $display("Passed the test case");
  end else $error("Failed. Outputs: %3d Expected Outputs: %3d", outputs, expected_outputs);

endtask

task wait_clocks(input integer num_clocks);
  #(num_clocks * CLK_PERIOD);
endtask
endmodule
